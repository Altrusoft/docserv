index.title = Välkommen till DocServ
index.services = Tillgängliga tjänster
index.service.version = returnerar versionsnummer för DocServe
index.service.templates = listar registrerade mallar
templates.registered = Registrerade mallar
